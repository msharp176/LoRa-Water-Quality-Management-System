** Profile: "SCHEMATIC1-rg_sweep"  [ C:\Users\mshar\Documents\capstone\simulation\Software-Defined Instrumentation Amplifier\Software_Defined_Instrumentation_Amplifier\Software_Defined_Instrumentation_Amplifier-PSpiceFiles\SCHEMATIC1\rg_sweep.sim ] 

** Creating circuit file "rg_sweep.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\cds_spb_home\cdssetup\OrCAD_PSpiceTIPSpice_Install\23.1.0\PSpice.ini file:
.lib "nom_pspti.lib" 
.lib "nom.lib" 

*Analysis directives: 
.DC LIN PARAM RG 1 100k 10 
.OPTIONS ADVCONV
.OPTIONS FILEMODELSEARCH
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
